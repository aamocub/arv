module arv (
    input wire logic clk_i,
    input wire logic rst_ni
);

endmodule
