// 
// ARV Core definitions.
//
// All parameters, types and functions used in the 'arv' core are defined here.

package arv_pkg;
    localparam integer unsigned PHY_ADDR_SIZE = 32;
    localparam integer unsigned VIRT_ADDR_SIZE = 64;
endpackage : arv_pkg
