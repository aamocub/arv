module arv #() ();
endmodule
