module tb_top;
    initial begin
        $display("Hello world\n");
    end
endmodule
