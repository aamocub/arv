// 
// RISC-V Specification definitions.
//
// All RISC-V related definitions should be defined in this package so that it can be easily
// included in all modules.

`ifndef RISCV_PKG_SV
`define RISCV_PKG_SV

package riscv_pkg;
    localparam integer XLEN = 32;
endpackage : riscv_pkg

`endif  // RISCV_PKG_SV
