module arv
    import arv_pkg::*;
    import riscv_pkg::*;
#(
) ();
endmodule
