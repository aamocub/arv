module arv_tb ();

endmodule
